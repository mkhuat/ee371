/*
Implements a simple Nios II system for the DE-series board.

Inputs: SW7−0 are parallel port inputs to the Nios II system
CLOCK_50 is the system clock
KEY0 is the active-low system reset
Outputs: LEDR7−0 are parallel port outputs from the Nios II system

*/
module Nios_processor (clk, reset, SW, LEDR, parallel_in, parallel_out, data_received, load, transmit_enable);
	
	// Inputs
	input clk;
	input [0:0] reset; // can assign this to KEY 0
	input [7:0] SW;
	input [7:0] parallel_in;
	
	// Outputs
	output [7:0] LEDR;
	output [7:0] parallel_out;
	output load, transmit_enable, data_received; 
	
	// Instantiate the Nios II system module generated by the Qsys tool:
	nios_sys u0 (
		.clk_clk                                    (clk),
		.leds_external_connection_export            (LEDR),
		.reset_reset_n                              (reset),
		.switches_external_connection_export        (SW),
		.load_external_connection_export            (load),
		.parallel_output_external_connection_export (parallel_out),
		.parallel_input_external_connection_export  (parallel_in),
		.data_received_external_connection_export   (data_received),
		.transmit_enable_external_connection_export (transmit_enable)  // transmit_enable_external_connection.export
	);

		
endmodule
