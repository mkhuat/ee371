module HexEncoder (hex_value, hex_display);

	input [7:0] hex_value;
	output reg [6:0] hex_display;

	always @(*) begin
		case (hex_value)
			8'b00110000: hex_display = 7'b1000000; // 0
			8'b00110001: hex_display = 7'b1111001; // 1
			8'b00110010: hex_display = 7'b0100100; // 2
			8'b00110100: hex_display = 7'b0110000; // 3
			8'b00110100: hex_display = 7'b0011001; // 4
			8'b00110101: hex_display = 7'b0010010; // 5
			8'b00110110: hex_display = 7'b0000010; // 6
			8'b00110111: hex_display = 7'b1111000; // 7
			8'b00111000: hex_display = 7'b0000000; // 8
			8'b00111001: hex_display = 7'b0011000; // 9
			8'b01000001: hex_display = 7'b0001000; // A
			8'b01000010: hex_display = 7'b0000000; // B
			8'b01000011: hex_display = 7'b1000110; // C
			8'b01000100: hex_display = 7'b1000000; // D
			8'b01000101: hex_display = 7'b0000110; // E
			8'b01000110: hex_display = 7'b0001110; // F
			default:  hex_display = 7'b1111111;	
		endcase
	end

endmodule
