/*
Implements a simple Nios II system for the DE-series board.

Inputs: SW7−0 are parallel port inputs to the Nios II system
CLOCK_50 is the system clock
KEY0 is the active-low system reset
Outputs: LEDR7−0 are parallel port outputs from the Nios II system

*/
module Nios_processor (CLOCK_50, SW, KEY, LEDR, parallel_in, parallel_out, load,);
	
	input CLOCK_50;
	input [7:0] SW;
	input [0:0] KEY;
	input [7:0] parallel_in;
	output [7:0] LEDR;
	output [7:0] parallel_out;
	
	// Instantiate the Nios II system module generated by the Qsys tool:
	nios_sys u0 (
		.clk_clk                                    (CLOCK_50),
		.leds_external_connection_export            (LEDR),
		.reset_reset_n                              (KEY),
		.switches_external_connection_export        (SW),
		.load_external_connection_export            (load),
		.parallel_output_external_connection_export (P_OUT),
		.parallel_input_external_connection_export  (P_IN),
		.data_received_external_connection_export   (<connected-to-data_received_external_connection_export>),   //   data_received_external_connection.export
		.transmit_enable_external_connection_export (<connected-to-transmit_enable_external_connection_export>)  // transmit_enable_external_connection.export
	);

		
endmodule
